module round();
endmodule;